`ifndef AXI_4_LITE_CONFIGURATION_V
`define AXI_4_LITE_CONFIGURATION_V

// Data bus details
`define C_AXI_DATA_WIDTH   32
`define C_REGISTERS_NUMBER 32

`endif